module CPU(tx, ty, tz, tula, acumulador, barramento, ulaout, entrada, clock);
	input wire clock;
	
	output [3:0] out;
	output [3:0] tx, ty, tz, tula, acumulador, barramento, ulaout, entrada;
	
endmodule
