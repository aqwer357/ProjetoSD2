module RegY(ulaout, acumulador, ty, clock);
	input wire clock;
	input wire [3:0] ulaout, ty;
	output reg [3:0] acumulador;
	
	parameter CLEAR = 4'd0;
	parameter LOAD = 4'd1;
	parameter HOLD = 4'd2;
	parameter SHIFTR = 4'd3;
	
	always@(posedge clock)
	begin
		case(ty)
			CLEAR: acumulador <= 4'd0;
			LOAD: acumulador <= ulaout;
			//HOLD: nada
			SHIFTR: acumulador <= acumulador >> 1;
		endcase;
	end
	
endmodule
